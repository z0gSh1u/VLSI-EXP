A SIMPLE CIRCUIT
.OPTIONS LIST NODE POST
.OP
.PRINT DC V(1) V(2) I(R1)
V1 1 0 DC=6V
R1 1 2 5
R2 2 0 10
.END